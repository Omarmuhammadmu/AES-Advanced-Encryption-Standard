package aes_package;
parameter BYTE = 8;
parameter WORD_SIZE = 32;
parameter DATA_WIDTH = 128;
parameter EXPANSIONED_KEY_SIZE = WORD_SIZE * 44;
parameter NUM_OF_ROUNDS = 10;

parameter MAT_NUM_ROW = 4;
parameter MAT_NUM_COLUMN = 4;
    
endpackage