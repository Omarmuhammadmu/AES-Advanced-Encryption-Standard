package aes_package;
parameter WORD_SIZE = 32;
parameter DATA_WIDTH = 128;
parameter EXPANSIONED_KEY_SIZE = WORD_SIZE * 44;
parameter NUM_OF_ROUNDS = 10;


// g operator typedef

// typedef union packed {
//     bit [WORD_SIZE-1:0] i_word;
//     bit [7:0] [3:0] byte_num;
// } wd_access;

    
endpackage