import aes_package::*;

module add_round_key (
    input  logic [DATA_WIDTH-1:0] data,
    input  logic [DATA_WIDTH-1:0] key,
    output logic [DATA_WIDTH-1:0] data_w_round_key 
);



endmodule